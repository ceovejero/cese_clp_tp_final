package param_package is

    constant    NUM_POINTS 		: integer := 4096;
	constant	MAX_AMPLITUDE 	: integer := 255;
	constant	ADDRES_BITS     : integer := 12;
	constant	AMPLITUDE_BITS  : integer := 12;

end param_package;

